------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : num32_play_sprite16x16.ppm 
--- Filas    : 512 
--- Columnas : 16 
--- Color    :  Blanco y negro. 2 niveles (1 bit)


-- 32 Imagenes, posiciones (5 bits mas significativos)
-- de 0x00 a 0x09: los numeros del 0 al 9
-- 0x0A: P
-- 0x0B: L
-- 0x0C: A
-- 0x0D: Y
-- 0x0E: S
-- 0x0F: T
-- 0x10: O
-- 0x11: W
-- 0x12: I
-- 0x13: N
-- 0x14: !
-- 0x15: :
-- 0x16: Mario
-- 0x17: Mario run
-- 0x18: Mario jump
-- 0x19: pacman
-- 0x1A: monster
-- 0x1B: monster afraid
-- 0x1C: cerezas
-- 0x1D: fresa
-- 0x1E: coche carreras hacia arriba
-- 0x1F: coche carreras diagonal


------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 16 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity memo_blue_16x16 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(9-1 downto 0);
    dout : out std_logic_vector(16-1 downto 0) 
  );
end memo_blue_16x16;


architecture BEHAVIORAL of memo_blue_16x16 is
  signal addr_int  : natural range 0 to 2**9-1;
  type memostruct is array (natural range<>) of std_logic_vector(16-1 downto 0);
  constant filaimg : memostruct := (
       "1111000000000111", -- 0x00 : 0
       "1110000000000011",
       "1100000000000001",
       "1100000110000001",
       "1100001110000001",
       "1100001110000001",
       "1100001100000001",
       "1100001100100001",
       "1100001000100001",
       "1100001001100001",
       "1100000001100001",
       "1100000011100001",
       "1100000011000001",
       "1100000000000001",
       "1110000000000011",
       "1111000000000111",
       "1111110000001111", -- 0x01 : 1
       "1111110000001111",
       "1111000000001111",
       "1111000000001111",
       "1100000000001111",
       "1100000000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011", -- 0x02 : 2
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1111111111000000",
       "1111111111000000",
       "1111000000000000",
       "1111000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000011111111",
       "1100000011111111",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011", -- 0x03 : 3
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1111111111000000",
       "1111111111000000",
       "1111110000000000",
       "1111110000000000",
       "1111110000000000",
       "1111110000000000",
       "1111111111000000",
       "1111111111000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1111000011111111", -- 0x04 : 4
       "1111000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111111111000000",
       "1111111111000000",
       "1111111111000000",
       "1111111111000000",
       "1100000000000000", -- 0x05 : 5
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000011111111",
       "1100000011111111",
       "1100000000000011",
       "1100000000000011",
       "1100000000000000",
       "1100000000000000",
       "1111111111000000",
       "1111111111000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1111000000000011", -- 0x06 : 6
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011111111",
       "1100000011111111",
       "1100000000000011",
       "1100000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1100000000000000", -- 0x07 : 7
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111111111000000",
       "1111111111000000",
       "1111111100000011",
       "1111111100000011",
       "1111111100000011",
       "1111111100000011",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111000000000011", -- 0x08 : 8
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1111000000000011",
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1111000000000011", -- 0x09 : 9
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000000",
       "1111000000000000",
       "1111111111000000",
       "1111111111000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1100000000000011", -- 0x0A : P
       "1100000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000011",
       "1100000000000011",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111", -- 0x0B : L
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111110000001111", -- 0x0C : A
       "1111110000001111",
       "1111000000000011",
       "1111000000000011",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000", -- 0x0D : Y
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111000000000011", -- 0x0E : S
       "1111000000000011",
       "1100000000000000",
       "1100000000000000",
       "1100000011111111",
       "1100000011111111",
       "1100000000000011",
       "1100000000000011",
       "1111000000000000",
       "1111000000000000",
       "1111111111000000",
       "1111111111000000",
       "1100000000000000",
       "1100000000000000",
       "1111000000000011",
       "1111000000000011",
       "1100000000000000", -- 0x0F : T
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111000000001111", -- 0x10 : O
       "1111000000001111",
       "1100000000000011",
       "1100000000000011",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "1100000000000011",
       "1100000000000011",
       "1111000000001111",
       "1111000000001111",
       "0000001111000000", -- 0x11 : W
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000000011000000",
       "0000000011000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "1100000000000011",
       "1100000000000011",
       "1111000000000011", -- 0x12 : I
       "1111000000000011",
       "1111000000000011",
       "1111000000000011",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111110000001111",
       "1111000000000011",
       "1111000000000011",
       "1111000000000011",
       "1111000000000011",
       "1100000011000000", -- 0x13 : N
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000000000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011000000",
       "1100000011111111", -- 0x14 : !
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1111111111111111",
       "1111111111111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1111111111111111", -- 0x15 : :
       "1111111111111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1100000011111111",
       "1111111111111111",
       "1111111111111111",
       "1111100000111111", -- 0x16 : Mario
       "1111000000000111",
       "1111000000011111",
       "1110000000000111",
       "1110000000000011",
       "1110000000000111",
       "1111100000000111",
       "1111110111111111",
       "1111110110111111",
       "1111110000111111",
       "1100101001010011",
       "1100000000000011",
       "1100000000000011",
       "1111000110001111",
       "1110001111000111",
       "1100001111000011",
       "1111100000110001", -- 0x17 : Mario run
       "1111000000000001",
       "1111000000011111",
       "1110000000000111",
       "1110000000000011",
       "1110000000000111",
       "1111100000001111",
       "1111110111011110",
       "0011111011101100",
       "0001111000010000",
       "1011010010000000",
       "1100000000000000",
       "1000000000011111",
       "1001111111111111",
       "1111111111111111",
       "1111111111111111",
       "1000111111110001", -- 0x18 : Mario Jump
       "1000100000010001",
       "1000000000000001",
       "1111000000001111",
       "1111000000001111",
       "1111100000001111",
       "1111100000011111",
       "1111100000011111",
       "1111100000011111",
       "0111110110111110",
       "0011110110111100",
       "0000110000110000",
       "0000001001000000",
       "0000000000000000",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111", -- 0x19 : Pacman
       "1111111111111111",
       "1111110000011111",
       "1111000000000111",
       "1110000100000011",
       "1110000000000011",
       "1100000000001111",
       "1100000001111111",
       "1100001111111111",
       "1100000001111111",
       "1100000000001111",
       "1110000000000011",
       "1110000000000011",
       "1111000000000111",
       "1111110000011111",
       "1111111111111111",
       "1111111111111111", -- 0x1A : Monster
       "1111110000111111",
       "1111000000001111",
       "1110000000000111",
       "1101100001100011",
       "1111110011110011",
       "1111110011110011",
       "1011110011110001",
       "1001100001100001",
       "1000000000000001",
       "1000000000000001",
       "1000000000000001",
       "1000000000000001",
       "1001000110001001",
       "1011100110011101",
       "1111111111111111",
       "1111111111111111", -- 0x1B : Monster afraid
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111",
       "1111110001001111", -- 0x1C : cherry
       "1111100000000011",
       "1111000111110001",
       "1110001111111000",
       "1111111111111100",
       "1111111111111101",
       "1110010111111111",
       "1100010010100111",
       "1000000100100011",
       "1000001000000001",
       "1001001000000001",
       "1000101001000001",
       "1100001000100001",
       "1110000100000011",
       "1111111110000111",
       "1111111111111111",
       "1111111111111111", -- 0x1D : Strawberry
       "1111000010000111",
       "1110000000000011",
       "1100000000000011",
       "1000000000000001",
       "1000000000000001",
       "1000000000000001",
       "1000000000000001",
       "1100000000000011",
       "1100000000000011",
       "1110000000000111",
       "1111000000000111",
       "1111100000001111",
       "1111110000011111",
       "1111111000111111",
       "1111111111111111",
       "1111111111111111", -- 0x1E : Racing car up
       "1111111111111111",
       "1111111111111111",
       "1111100000011111",
       "1111100000011111",
       "1111111001111111",
       "1111111001111111",
       "1111110000111111",
       "1111110000111111",
       "1111100000011111",
       "1111100000011111",
       "1111000000001111",
       "1111000000001111",
       "1111100000011111",
       "1111111111111111",
       "1111111111111111",
       "1111111111111111", -- 0x1F : Racing car diagonal
       "1111111111111111",
       "1111111111011111",
       "1111111110001111",
       "1111111110000111",
       "1111111110000011",
       "1111111100000111",
       "1111110000111111",
       "1110000001111111",
       "1100000001111111",
       "1100000011111111",
       "1110000011111111",
       "1111000001111111",
       "1111100011111111",
       "1111111111111111",
       "1111111111111111"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
   end if;
  end process;

end BEHAVIORAL;
